//`define ISE
`define SIMULATION

`ifdef ISE
`define ISE_OR_SIMULATION
`endif

`ifdef SIMULATION
`define ISE_OR_SIMULATION
`endif


