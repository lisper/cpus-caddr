`define ISE
//`define ISE_OR_SIMULATION
