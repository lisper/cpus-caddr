//

module mmc_disk(
		input mmc_cs, input mmc_di, output mmc_do, input mmc_sclk
		  );
   
endmodule // mmc_disk
